`timescale 1ns / 1ps

module integrationConv_TB ();

    // === 参数配置 ===
    parameter DATA_WIDTH = 16;
    parameter ImgInW = 32;
    parameter ImgInH = 32;
    parameter DepthC1 = 6;
    parameter Conv1Out = 32;
    parameter Conv1Kernel = 5;
    parameter MvgP1out = 16;
    parameter DepthC2 = 16;
    parameter Conv2Out = 12;
    parameter Conv2Kernel = 5;
    parameter MvgP2out = 6;
    parameter DepthC3 = 32;
    parameter Conv3Out = 6;
    parameter Conv3Kernel = 3;
    parameter MvgP3out = 3;

    // === 信号定义 ===
    reg clk, reset;
    reg  [                          ImgInW*ImgInH*DATA_WIDTH-1:0] CNNinput;
    reg  [      1*Conv1Kernel*Conv1Kernel*DepthC1*DATA_WIDTH-1:0] memory1     [ 0:6-1];
    reg  [      1*Conv1Kernel*Conv1Kernel*DepthC1*DATA_WIDTH-1:0] Conv1F;
    reg  [DepthC1*Conv2Kernel*Conv2Kernel*DepthC2*DATA_WIDTH-1:0] memory2     [0:16-1];
    reg  [DepthC1*Conv2Kernel*Conv2Kernel*DepthC2*DATA_WIDTH-1:0] Conv2F;
    reg  [DepthC2*Conv3Kernel*Conv3Kernel*DepthC3*DATA_WIDTH-1:0] memory3     [0:32-1];
    reg  [DepthC2*Conv3Kernel*Conv3Kernel*DepthC3*DATA_WIDTH-1:0] Conv3F;
    wire [              MvgP3out*MvgP3out*DepthC3*DATA_WIDTH-1:0] iConvOutput;

    integer i, fd, code;

    // === DUT 实例化 ===
    integrationConv uut (
        .clk        (clk),
        .reset      (reset),
        .CNNinput   (CNNinput),
        .Conv1F     (Conv1F),
        .Conv2F     (Conv2F),
        .Conv3F     (Conv3F),
        .iConvOutput(iConvOutput)
    );

    localparam PERIOD = 10;
    // === 时钟产生 ===
    initial clk = 0;
    always #5 clk = ~clk;  // 100MHz 时钟

    // === 仿真控制 ===
    initial begin
        $display("==== Start Simulation ====");
        reset = 1;
        CNNinput = 0;
        Conv1F = 0;
        Conv2F = 0;
        Conv3F = 0;

        // 保持复位
        #20;
        reset = 0;

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv1_hex.txt", "r");
        for (i = 0; i < 6; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory1[i]);
        end
        for (i = 0; i < 6; i = i + 1) begin
            Conv1F[i*5*5*16+:5*5*16] <= memory1[DepthC1-1-i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv2_hex.txt", "r");
        for (i = 0; i < 16; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory2[i]);
        end
        for (i = 0; i < 16; i = i + 1) begin
            Conv2F[i*5*5*6*16+:5*5*6*16] <= memory2[DepthC2-1-i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv3_hex.txt", "r");
        for (i = 0; i < 32; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory3[i]);
        end
        for (i = 0; i < 32; i = i + 1) begin
            Conv3F[i*3*3*16*16+:3*3*16*16] = memory3[DepthC3-1-i];
        end

        CNNinput = 16384'h33883525368736f735e633272f472c04298628042a872c852d862e87300431a633a834e53586358634d534743404324630642ec72ec730e534143606377737673676370737a837d83727351531652c4425052004200424042505260629052c442f47314533273454341434443505359634e5332730e52f472f88310532a73414377737983777379837e83788359631862a87240422062606270724042004240428852c442fc8326634443575367636c7368736c736d7362634c531a62f072e4636d73656366636f737c8385c3854369733882ec72a062707240420041c041c04200427072cc530c5342435e6363634e53307342435653666371736b735d634f536c736763717381c386c387438b5388d3788355532e72fc82b88288525052206240428852d053186350536b73697347430642e062f073165348536c7380c380437c8385c387c38b538fd38d538a538ad38b53864379835a633e831e630c52fc83004302430e533e8365637a837a836a73505338831e6318632c73535372737f8388d390538d53874383c37c83798384438d538fd38dd3854379836d7363635b635e63616363636d737f8384c383437c837073505324630a531e634a536873767390d391d388536d73485324632e735653788386438d538bd388d3874386c3834385c388d388d388538a538a5386c380c371734442f472a062c043044347435f6395d3925383c354530442b882c042f8832e735a6381438b538cd38c538d538ad389538ad38dd38c538dd387c381c37e8371734c531c62f472c042986306434443975396538c5363630852a0629052b072dc631e63616384c38c538cd38ed38d53895389538a5383437983656353534d5354535453555351533e8310531e63474399e39ce392d37c834c530042c442cc52e873125352537c8389538dd392d391538d538dd387435d6334731252fc82e873044320634743616371736c7369736b7399e39ae3965390d38543565338833a8347434d53626380c38b538ed38ed38ed38f538cd37a833a82ec72c042986280429862cc5304433883646381c3854380c397d394d394d3986396538a53824380c3814380c3834387438ad388d3814382438a53874363631a62cc5290526062206240428042a062dc6328735c6377737b8392d38c538d5390538ed38a5384c3834382c382c38743885386c380c37073737385c388536c732462c442707240420042004240427072b072fc8345436b7377738d53834376736a735f635a63525355535863575364636c73747375736e73757388538fd380c33a82d05260622062004200425052b8830243367359637173757382c3606342431e630e53105316531a631653165328733e834c5352535553676385c38f5383434c52f472804200422062b073024338835a6370737d837f83727368733072f472d452c442c042d052d452d052e062f8830c531a6322632e734b53737385c382c36a7343430a52e0630243434362637773844389538a53864377735e631a62c442804260624042707270728042a062c442d452f07306430e533a83687384c389d3885380c371736c73757381c3864388538743854389d388d382c37b834c52ec724041c0420042004200420042404260628852c442e8730c534853757388d38cd390d39253935393d393538fd38e538ed38a53814385c3895388d37c83747354531e62cc5220600000000000000002004200427072e4633473656384438853844387438f5392d3935393d39553965394538e5388d387438a538bd35b636c7380437e835f633272fc82c4429052707250527072b073044349537883895387437f8382438bd390d390538e538d538bd3895386c384c381c388d38e5363635d63707381c382c380436f7364635453367326633e8344434c536c7385c38cd38bd3885387c385c3824376736163515349534a534e5351535753717384436c73505340434043485359637573864387c380c37c838143824383c38b538b538ad38b5388d37b8359633e831862f882e062cc52cc52d862e8730443206343436f734c530a52b882a872d053186343435d637883844387c389d38bd38e538b538b5388d3798349530a52d052b0729862707250524042606280429862a872d0537f836873454304429052404250528852cc531c635a6376737f838143854386c38b5386435f630a52a062a062a87288524042206220622062505240426062c0437273788373735d633672f882c852905260629862f47328734c53626372737b83874386c36a733072d862a87298627072004200420042206250528852d8631e63495367637983804378835a63464332731c630442b882a8730243424365637b8386438bd38b537d8346430a52d862a0628852a062e0630243004322634d53697310534b536f738343854382437f837b83747364634b53404332733a835863788382c38543895387c37a836c7358634143434346435963697365636b737273747322634c536b7381c3874388538a5389d388d38a538d538b5382c37173687373737a837b837983767372737473717365635d63565354535653586356534e53485359636d737b8382c3874388d385c378836c7372737f8385c389d387c380c37c83788377737373636346432c731a630642ec72e062d452d052e062f472f072e8737e83824385438643874386c373734a53165300430a53206340434853434343434743535361635f6343430c52c8526062505250522062004240428042885280438bd3895386c385c3854383c36f734342f472b882a87298628852804280428852a872e46322634b53505344431a62d45288524041c041c041c04200422062206;

        // 运行一段时间
        #(75050 * PERIOD);

        $display("==== Simulation Done ====");
        $display("[%0t] iConvOutput = %h", $time, iConvOutput);
        $stop;
    end

endmodule
