// CNN_FGPA\CNN_FPGA.sim\sources_1\new\convLayerMulti.v
`timescale 1 ns / 1 ps

module convLayerMulti_TB();

parameter DATA_WIDTH = 16;
parameter D = 1;  //Depth of image and filter
parameter H = 32;  //Height of image
parameter W = 32;  //Width of image
parameter F = 5;  //Size of filter
parameter K = 6;  //Number of filters applied
parameter P = 0;  //Number of padding pixels

reg clk, reset;
reg [0:D*H*W*DATA_WIDTH-1] image;
reg [0:K*D*F*F*DATA_WIDTH-1] filters;
wire [0:K*(H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH-1] outputConv;

localparam PERIOD = 4;

integer i,j,k;

always
	#(PERIOD/2) clk = ~clk;

convLayerMulti #(
    .DATA_WIDTH(DATA_WIDTH),
    .D(D),
    .H(H),
    .W(W),
    .F(F),
    .K(K),
    .P(P)
)
UUT 
(
	.clk(clk),
	.reset(reset),
	.image(image),
	.filters(filters),
	.outputConv(outputConv)
);
	
initial begin 
	#0
	clk = 1'b0;
	reset = 1'b1;
	#1
	reset = 1'b0;
	// input image = 1*32*32*16 = 16384 bit
	// expected output = 6*32*32*16 = 98304 bit
	 image = 16384'h56ae58d657fd5b2a58565bde56b73c08535f59044a835bcd59525be24d6f5086570559f55b0f593d555e4b5b5bdb375348d45b52561a51675049599353195b0b554b512b3cd64d0358ff45eb5b2b55e75ab14dd855305acc554b5b2f3d6250b656be5470562f556d5a955ab154f953bf5b4a543055fe592b5a81599b503a554858a859055440561c4c00460f54945a595a334e00557a5bdd582c4fbf526e565b5a9d59d55b8e5bb459a74f7c5b3857ea5a81504558c64e423d5658c359ed5ba14a124e9a561d5ba04d4f576b54795a9455e45a96597c58fa573f5b505a3859415a215a325b825aff580a5815594a572c5abf5bf659fc588a5b9b58f550294bd5575b4dc758a45b265afe5abe577054e95acb529b585f59ae4df155f44cbc58df580159c05932597c4cbc532d5ae658e3511956c95678508e5548597f532f506853265a0758a84a8e5860588f55e158a55ab65bb83a284d4458e859c054e4561a50d94208570e5bc1495f4d1f5b3d5acf598055d35741589550ad541e48705a9a5b054d395a8158025a5d5be1597756635bbb58f155205a6759635685594b569356495b005aad543e4ee94a18582e544558d458ff55cd4bd85946584f53e159b8531d45e6580956e85b07592e5ba75a0657a754ca5b005a1458f553e24d8751e1599f5ad1514350e65194596850365b4c5573534d55885b6454dd46b953d55b625a905aee5506558f57ba4d875ae3546c5b7c5a71546a5537587f58db544647524edb5ada52144d855a89599455df5abc57f653c154ba4d9755e0565e5b5959b759b9540b52ec543952565a5742524f54562c365a5a415a1159f65b595a845b534572580949205b445bcd516954b057fa5aa05820587947b759ef576f58b15bb8542c54b65947523c49fd552f4c815b9b59f9584e541c5acc547954ff5b6c54645a5634405b314e8d54d1531357cf5a3b4c08544e50055b3c545758ac52b959134869543e57de5b385a9f55f55a0f50a758df5b415709502e4dec54da5af85ac655c55b7055b559055a6b5a145ab35ac159c3551d5018560a575c58655473587759d645ef5a2e50345a9458e05a0a4993440257325bf759365b725992566559264b6f58355a6758085a4a4d564ba64c1558235b1f5a8b4daa5a9a551c54fa54e4485f580a567c53775b4f5a414b7e57fa4e36539f549e59795a095a435834566353ae5aea54a156a35951592c5b995723589f5610578b46a651f34dba58e356f257f44c2255f3580f5be352cd5b9c4d545abe54e54cdf58d1517c576359da560659f5583054755a2759604965587a5964583b57074b25480e563f5bce57eb590e5b3a4fb65a2c57de5a495b1d5be25acc58fe50b25b2a5947562758d45b2f59d45a4350bc5b3b595c5b4d5b305447583a4b435b6d5a4258c147fe59fc581d5131583b5b5c5910584d594151065be154f85615584f50975b41583656e94b13581c58894fd34f2045b654885b7158a657f658585a8c5a245af85513595d36cc455a3a08599e4e0c55605b6653cd42825a525b0f5b8e5b29591e591359fe592a536d57c24fd6596e54e45af45bb05acd50e65aea5507583b57ca5acf5b6b592b5af159df5888579c5a1056ff59d2583a584555db59b45084546143404c9b5811591b54755b0e3a9150174c2f5ad155ba492f5ac25b875640575f48e859d05ad05bef59ed43bd5b154dd558605a7a545c5a115880569157e059c7552f588f58005a5157f35ac85be958f8500259624b394c8f594751865a01457140155bc558fa5796366b4e0755894d195a0752d255fd5a0150b759ef42f55a5e5866599b5bbc541c5bc559fd59f754135afb4da75b4255055bad540d55e25b1a460258274ffd4f1e54ba5a695b3f5901593c5bdf58f35b065b195557579154c456db5ade4947550d5ac15bd05bd4562c5ae3598f5a545b875b4e5b3451c65ae358224d375a4a5484589d56e34b40593444c35b3053d955a357a159725a0048a55b0b588956485a8259b65a4654e85acc5b605305565a587654795558552255f14d8d55ff55ba5af15af456265a604d0250d154ad5474517a585c55cc54f959f957f94f304d07594d4f6a5ad35bf85694574c523a58e957d75b8b57f95bef5b9b52d24adc56015a1a5900586959a452b759f755dd573e513d53d356de59ad59bd58fb549b5b7b543d5b8e55e8572958cf59d85bd059665a8357735a335bef517b54fa595a5b8c57a3581d4dfb59c35b9f5246566458c5526651a3575c556b570f5944582e56dd560159ac57df4d535b785b025780545058565b1f5aa1598b526958e5506657d95b0259c05b55566159eb56f853ed5a8a59515ae252b3516e4d7b4ed156d34d0d52355a8a55e9546356e9594a5985508f490f58933c545ba1526d59265b16521c553e571c5b3050de5b5d5afb57f6488552225a5757ba575f580555a158b758005844573c53cf5a5a59a559025a804b7450c354a058f759cd502f5a8555ac58aa5a3358a056b353e44e0c51d2585e597757ee50b65709575558c1589a50ac5ae8581e57ce5422513c4cf45a2f52bc594e5b0d53e05a5355f7542d4cbc5ad555275a9b5a67590054cc58ed50fe59b4542d554d557e5a6d586c59385b2e58c759b150935a4a597752ec55f2597e486859b65a82545454915bb62ed559a45b115366591351b453b959bd56f75a71512c563653bc5a69565d59fd54dd59c85b3e5a3e520c514a59ac59785aef3a2b5ac356fa574e5a7d546254a95933590a59eb5150582156bf5b665a36560b5a705be659405a0a59f95be25bf04d9f581e55985927591b4d1f580858a35aea565458ac5b43559656d452365a9d5ad2491858da5a465847;
     // filters = 6*1*5*5*16 = 2400 bit
	 filters[0*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'ha48c311e37d231da336d374fb2e7b18e318ab2c8b52a378cae7bb107b3f2b72820c4b698b706b2baa0a6b4af349935adb59a;
  	 filters[1*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h34c1b654369c31a2b79836203188b58435f536722868b4e6b12b3441b6b3369fae129c8b337ca97934f131fc33742147379d;
	 filters[2*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'hb0ae200c330eb6353004b6373771b4ea35f29f1333afb42c2d61b2d12da633afb503b580277634f9b54db62e36e834d7b5af;
	 filters[3*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'hb50734932eb12b24b56faeafb5f3375728acb6df3773300a347f350c2f1a2c409b5234a235d4307eb5b59727366d33fdaec4;
	 filters[4*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'hb206a509ae5a2f3aaf48b0ffafa7359f2b5a34e436cf3459345b369fb477b66e3438b3e4a0043072ac50237731f32a61378b;
	 filters[5*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h326734f92d43b665afd837d6b45c30bb331bb2a123112e28b621b061b54bb45cb681242bb6093699353fb7dc343a327d376e;
	#(PERIOD)

	// reset = 0;
	
	#(3*1793*PERIOD)
	// Display output
    for (k = 0; k < 6; k = k + 1) begin
        $display("Kernel %d result is %h ", k+1, outputConv[k*(H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH +: (H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH]);
        $display("\n");
    end
	$stop;
end

endmodule
