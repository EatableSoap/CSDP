// CNN_FGPA\CNN_FPGA.sim\sources_1\new\IntegrationConvPart.v
// `timescale 100 ns / 10 ps

module IntegrationConvPart_TB ();
endmodule