// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\MaxPoolSingle.v
`timescale 1 ns / 10 ps

module MaxPoolSingle_TB ();

    parameter DATA_WIDTH = 16;
    parameter InputH = 28;
    parameter InputW = 28;
    parameter Depth = 1;

    reg     [        InputH*InputW*Depth*DATA_WIDTH-1:0] aPoolIn;
    wire    [(InputH/2)*(InputW/2)*Depth*DATA_WIDTH-1:0] aPoolOut;
    integer                                              i;

    MaxPoolSingle #(
        .DATA_WIDTH(DATA_WIDTH),
        .InputH(InputH),
        .InputW(InputW),
        .Depth(Depth)
    ) UUT (
        .aPoolIn (aPoolIn),
        .aPoolOut(aPoolOut)
    );

    initial begin
        #0
        // aPoolIn = 28*28*1*16 = 12544 bits
        aPoolIn = 12544'h4000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004000440040004400400044004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200450042004500420045004200;

        #10
        // $displayh(outMaxPool[i*16+:16]);
        $display(
            "Result (hex): %h", aPoolOut[i*16+:16]
        );
        $stop;
    end

endmodule
