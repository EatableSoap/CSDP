// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\activationFunction.v
//`timescale 100 ns / 10 ps

module activationFunction_TB ();

parameter DATA_WIDTH = 32;
parameter OUTPUT_NODES = 32;

reg clk, reset, en;
reg [DATA_WIDTH*OUTPUT_NODES-1:0] input_fc;
wire [DATA_WIDTH*OUTPUT_NODES-1:0] output_fc;


localparam PERIOD = 100;

always
    #(PERIOD/2) clk = ~clk;

activationFunction #(
    .DATA_WIDTH(DATA_WIDTH),
    .OUTPUT_NODES(OUTPUT_NODES)
)
UUT
(
	.clk(clk),
	.reset(reset),
	.en(en),
	.input_fc(input_fc),
	.output_fc(output_fc)
);

initial begin
	#0
	clk = 1'b0;
	reset = 1'b1;
	en = 0;
    // input: 32*32 = 1024 bit
	input_fc = 1024'b1000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000;

	#PERIOD
	reset = 0;
	en = 1'b1;

	#PERIOD
    // input: 32*32 = 1024 bit
	input_fc = 1024'b0100000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000;

	#PERIOD
	$stop;
end

endmodule