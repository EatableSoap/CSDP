// CNN_FGPA\CNN_FPGA.sim\sources_1\new\Lenet.v
`timescale 1 ns / 1 ns

module Lenet_TB ();

    reg [32*32*16-1:0] input_ANN;

    reg clk, reset;
    wire    [             3:0] output_ANN;
    reg     [    5*5*6*16-1:0] Conv1F;
    reg     [         400-1:0] memory1    [ 0:6-1];
    reg     [ 5*5*6*16*16-1:0] Conv2F;
    reg     [    5*5*6*16-1:0] memory2    [0:16-1];
    reg     [3*3*16*32*16-1:0] Conv3F;
    reg     [   3*3*16*16-1:0] memory3    [0:32-1];

    integer                    i;
    integer                    code;
    integer                    status;
    integer                    fd;

    localparam PERIOD = 4;

    always #(PERIOD / 2) clk = ~clk;

    initial begin

        #0 clk = 1'b0;
        reset = 1'b1;

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv1_hex.txt", "r");
        for (i = 0; i < 6; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory1[i]);
        end
        for (i = 0; i < 6; i = i + 1) begin
            Conv1F[i*5*5*16+:5*5*16] <= memory1[5-i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv2_hex.txt", "r");
        for (i = 0; i < 16; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory2[i]);
        end
        for (i = 0; i < 16; i = i + 1) begin
            Conv2F[i*5*5*6*16+:5*5*6*16] <= memory2[15-i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv3_hex.txt", "r");
        for (i = 0; i < 32; i = i + 1) begin
            code <= $fscanf(fd, "%h", memory3[i]);
        end
        for (i = 0; i < 32; i = i + 1) begin
            Conv3F[i*3*3*16*16+:3*3*16*16] = memory3[31-i];
        end


        // label:0
        // #(PERIOD / 2) reset = 1'b0;
        // input_ANN = 16384'h33883525368736f735e633272f472c04298628042a872c852d862e87300431a633a834e53586358634d534743404324630642ec72ec730e534143606377737673676370737a837d83727351531652c4425052004200424042505260629052c442f47314533273454341434443505359634e5332730e52f472f88310532a73414377737983777379837e83788359631862a87240422062606270724042004240428852c442fc8326634443575367636c7368736c736d7362634c531a62f072e4636d73656366636f737c8385c3854369733882ec72a062707240420041c041c04200427072cc530c5342435e6363634e53307342435653666371736b735d634f536c736763717381c386c387438b5388d3788355532e72fc82b88288525052206240428852d053186350536b73697347430642e062f073165348536c7380c380437c8385c387c38b538fd38d538a538ad38b53864379835a633e831e630c52fc83004302430e533e8365637a837a836a73505338831e6318632c73535372737f8388d390538d53874383c37c83798384438d538fd38dd3854379836d7363635b635e63616363636d737f8384c383437c837073505324630a531e634a536873767390d391d388536d73485324632e735653788386438d538bd388d3874386c3834385c388d388d388538a538a5386c380c371734442f472a062c043044347435f6395d3925383c354530442b882c042f8832e735a6381438b538cd38c538d538ad389538ad38dd38c538dd387c381c37e8371734c531c62f472c042986306434443975396538c5363630852a0629052b072dc631e63616384c38c538cd38ed38d53895389538a5383437983656353534d5354535453555351533e8310531e63474399e39ce392d37c834c530042c442cc52e873125352537c8389538dd392d391538d538dd387435d6334731252fc82e873044320634743616371736c7369736b7399e39ae3965390d38543565338833a8347434d53626380c38b538ed38ed38ed38f538cd37a833a82ec72c042986280429862cc5304433883646381c3854380c397d394d394d3986396538a53824380c3814380c3834387438ad388d3814382438a53874363631a62cc5290526062206240428042a062dc6328735c6377737b8392d38c538d5390538ed38a5384c3834382c382c38743885386c380c37073737385c388536c732462c442707240420042004240427072b072fc8345436b7377738d53834376736a735f635a63525355535863575364636c73747375736e73757388538fd380c33a82d05260622062004200425052b8830243367359637173757382c3606342431e630e53105316531a631653165328733e834c5352535553676385c38f5383434c52f472804200422062b073024338835a6370737d837f83727368733072f472d452c442c042d052d452d052e062f8830c531a6322632e734b53737385c382c36a7343430a52e0630243434362637773844389538a53864377735e631a62c442804260624042707270728042a062c442d452f07306430e533a83687384c389d3885380c371736c73757381c3864388538743854389d388d382c37b834c52ec724041c0420042004200420042404260628852c442e8730c534853757388d38cd390d39253935393d393538fd38e538ed38a53814385c3895388d37c83747354531e62cc5220600000000000000002004200427072e4633473656384438853844387438f5392d3935393d39553965394538e5388d387438a538bd35b636c7380437e835f633272fc82c4429052707250527072b073044349537883895387437f8382438bd390d390538e538d538bd3895386c384c381c388d38e5363635d63707381c382c380436f7364635453367326633e8344434c536c7385c38cd38bd3885387c385c3824376736163515349534a534e5351535753717384436c73505340434043485359637573864387c380c37c838143824383c38b538b538ad38b5388d37b8359633e831862f882e062cc52cc52d862e8730443206343436f734c530a52b882a872d053186343435d637883844387c389d38bd38e538b538b5388d3798349530a52d052b0729862707250524042606280429862a872d0537f836873454304429052404250528852cc531c635a6376737f838143854386c38b5386435f630a52a062a062a87288524042206220622062505240426062c0437273788373735d633672f882c852905260629862f47328734c53626372737b83874386c36a733072d862a87298627072004200420042206250528852d8631e63495367637983804378835a63464332731c630442b882a8730243424365637b8386438bd38b537d8346430a52d862a0628852a062e0630243004322634d53697310534b536f738343854382437f837b83747364634b53404332733a835863788382c38543895387c37a836c7358634143434346435963697365636b737273747322634c536b7381c3874388538a5389d388d38a538d538b5382c37173687373737a837b837983767372737473717365635d63565354535653586356534e53485359636d737b8382c3874388d385c378836c7372737f8385c389d387c380c37c83788377737373636346432c731a630642ec72e062d452d052e062f472f072e8737e83824385438643874386c373734a53165300430a53206340434853434343434743535361635f6343430c52c8526062505250522062004240428042885280438bd3895386c385c3854383c36f734342f472b882a87298628852804280428852a872e46322634b53505344431a62d45288524041c041c041c04200422062206;
        
        //label:6
        // input_ANN = 16384'h30042fc8302430a530852fc82f072e872e872d052c042a872b0729052a06298629862a062c442dc6310533e8379838a537d83747367634f5326631a6332735252ec7300430a52f882e062e462e062e062dc62c852c852c442c442b882b882986290529862b882cc52e0630e5338833473404340432a731e630e531e63327336730443024304430242f47300430442fc82e872dc62e462dc62d862c442b072b072c442c442c442c042c852e062ec72fc8312530c5308530c530a531453145306430242f882e462ec72f072fc830042ec72e462e872e872e062d452c042b072cc52e062e062c042a872b882c852d862ec72f882f472f47308530e5318632c733882f472f472e872f4730042f072e462e062dc62dc62dc62d452c852c042c442dc62e872d452a872b072c442cc52e462f472ec730443064306431453145318632662f072f472f072f072fc82ec72d862d862d862dc62d452d452e872e062d452cc52c042a06290529862b882cc52d862e872f472fc82f073004314531053064304430042f8830242fc82f882f882e872d452d452e062e062d452c852c442cc52cc52b07298628852a872b072c042cc52e062ec72f882e062e462f072f882fc830442e872f4730042e872f072f882f072d862d862e462ec72dc62cc52c852d862d452b882b882b072b072b072c852d052e462ec72f072fc83085304430c5314530852fc82e872f882f073004308530042ec72ec72ec72ec72f882e462d052cc52b882b882a8729862a872b072c042c852dc62e062dc62f88334733c831253004300430443105308530c531e6332732e7322631a631253085302430042f472f472cc52c442c042b072b882b882b882b882c852d862dc62e87308532263165308530c531a633e83545372738443824376736e7370737883687353534143226310530642e872d052c042b882c042b882b882cc52d862e062ec7312531c63085304430e5336736f7389d38cd394d395d393d39253975397d393d38cd37173495328732c731862ec72c852b072b882c442c852e872fc82f472e462ec7302430643085320635a6383c38cd3925397d395d396d39963935389d38ad38b5388d381c36a7350533a830e52dc62c852d05300432063464334730042d862e462f073085310533a83206348536b7387c38e5390d38e538cd38c539253965394d390538fd390d38dd377734c533273145304432a73596356533882f472e062f072f072e462f8832262f07320633e833c8346435c6357534e5368736763687369737b838dd391538c5386c381c373735c6344434853525340430042e872ec72ec72f073004300430042fc82f072e872f88310530a530c5322632663186308531e635c63757381438a5391d38d538c5380c35b6345433c831252f88306430242f472f4730c5310530852fc82fc82f472f882f072e062f072fc82f882f882f883064322633e83525366636b73767386c371735a633e830852dc62e0630242fc830e53145328732e731e6300430852fc82e872f472f882f882e872dc62f07304430242fc83024308531c6338835b636973737357532c730852dc62cc52d452e873004310530c53226324630642fc82e462e872e872f8830642fc82e8730042fc82dc62e462d862e062f0730443125326633673414344431252dc62d052e463064310530a5300430c5316531a62f882ec72f472fc8300430242f072dc62e062ec72e872d052d452dc62dc62dc62d862e46316535e635c632a7308530042e462e06302430a52f882fc830e5357531e63024306430e530a52f472ec72f472e462dc62e062d052d452d452cc52dc62e872e0631c63636367634f533473347328731e632663327322630242f0735c632a7302430a530c52fc82f072f8830642f072d452d052d452dc62d452d862dc62e062e06310534b5363636563656364636d7371736b735c634c531862dc634743145308530a530242f883064324633e8332730c530242f072e062d452e872f882f882e063105343434d536d737b837e838043804380437e836e73596332730a52f882f472ec72ec72e872e4630c532e7330730e530e5318631e62f882d052d862d862d052d86312534853666371737273757381c38c5390538e538bd37f82e872e462dc62d862d052e462e062d452e462e462ec72f8830e5324630c52e872e062e062d052b882f0732c733673464352535f636a7382438fd392d393538e52dc62d862d052d862e062e872f882f072d862d452e872f072e872e062e872f47304430852dc62c042d862f4730c53105318632c733a834b535353666384c38dd2e062e462dc62ec72f472e872e462e462e872cc52d052e062dc62e872fc82f073004314530242c442a872c442dc62e062f072e062f47300430043347352536562dc62e062f072f8830643125314531a630a52ec72d862d052d452dc62dc62f472f47300430c52ec72cc52c042b882d452d452d452d862dc62f883004322635352d052d052d862f0730c53347354536463515334730a52d862c042c442cc52cc52d052f8830a52e462c852b882c442d452e062dc62e062dc62e462f07306433672d862d862f07318634d536d7380c3885385c36a7345430c52c852c442cc52d052c852d452c852c442c042c042d862e462e462e062e872e462e462dc62f4731452d45300433473636382c385c385c38b5386436a732c72e462c852c042b882b882cc52cc52b882a872b882c442d052d862dc62e062ec72e462e872e872f473044300433883606377737d8383c387c3814361633e82fc82c852c852c852d452cc52cc52d452c442b882c442b882c852d862dc62dc62e872f47304430852fc83004;
        // #((75050 + 20 + 550) * PERIOD);
        // #(PERIOD * 100);

        fd = $fopen("D:/Material/CSDP/Data/small_test_image.txt", "r");
        for (i = 0; i < 10000; i = i + 1) begin
            #(PERIOD / 2) reset = 1'b0;
            #(PERIOD / 2);
            status = $fscanf(fd, "%h", input_ANN);
            #((75050 + 20 + 550) * PERIOD) #(PERIOD * 100) #(PERIOD / 2) reset = 1'b1;
            #(PERIOD / 2);
        end

        $stop;

    end

    Lenet UUT (
        .clk        (clk),
        .reset      (reset),
        .CNNinput   (input_ANN),
        .Conv1F     (Conv1F),
        .Conv2F     (Conv2F),
        .Conv3F     (Conv3F),
        .LeNetoutput(output_ANN)
    );

endmodule
