// CNN_FGPA\CNN_FPGA.sim\sources_1\new\Lenet.v
`timescale 1 ns / 1 ns

module Lenet_TB ();

    reg [32*32*16-1:0] input_ANN;

    reg clk, reset;
    wire    [             3:0] output_ANN;
    reg     [    5*5*6*16-1:0] Conv1F;
    reg     [         400-1:0] memory1    [ 0:6-1];
    reg     [ 5*5*6*16*16-1:0] Conv2F;
    reg     [    5*5*6*16-1:0] memory2    [0:16-1];
    reg     [3*3*16*32*16-1:0] Conv3F;
    reg     [   3*3*16*16-1:0] memory3    [0:32-1];

    integer                    i;
    integer                    code;
    integer                    status;
    integer                    fd;

    localparam PERIOD = 4;

    always #(PERIOD / 2) clk = ~clk;

    initial begin

        #0 clk = 1'b0;
        reset = 1'b1;

        // label:0
        // input_ANN = 16384'h33883525368736f735e633272f472c04298628042a872c852d862e87300431a633a834e53586358634d534743404324630642ec72ec730e534143606377737673676370737a837d83727351531652c4425052004200424042505260629052c442f47314533273454341434443505359634e5332730e52f472f88310532a73414377737983777379837e83788359631862a87240422062606270724042004240428852c442fc8326634443575367636c7368736c736d7362634c531a62f072e4636d73656366636f737c8385c3854369733882ec72a062707240420041c041c04200427072cc530c5342435e6363634e53307342435653666371736b735d634f536c736763717381c386c387438b5388d3788355532e72fc82b88288525052206240428852d053186350536b73697347430642e062f073165348536c7380c380437c8385c387c38b538fd38d538a538ad38b53864379835a633e831e630c52fc83004302430e533e8365637a837a836a73505338831e6318632c73535372737f8388d390538d53874383c37c83798384438d538fd38dd3854379836d7363635b635e63616363636d737f8384c383437c837073505324630a531e634a536873767390d391d388536d73485324632e735653788386438d538bd388d3874386c3834385c388d388d388538a538a5386c380c371734442f472a062c043044347435f6395d3925383c354530442b882c042f8832e735a6381438b538cd38c538d538ad389538ad38dd38c538dd387c381c37e8371734c531c62f472c042986306434443975396538c5363630852a0629052b072dc631e63616384c38c538cd38ed38d53895389538a5383437983656353534d5354535453555351533e8310531e63474399e39ce392d37c834c530042c442cc52e873125352537c8389538dd392d391538d538dd387435d6334731252fc82e873044320634743616371736c7369736b7399e39ae3965390d38543565338833a8347434d53626380c38b538ed38ed38ed38f538cd37a833a82ec72c042986280429862cc5304433883646381c3854380c397d394d394d3986396538a53824380c3814380c3834387438ad388d3814382438a53874363631a62cc5290526062206240428042a062dc6328735c6377737b8392d38c538d5390538ed38a5384c3834382c382c38743885386c380c37073737385c388536c732462c442707240420042004240427072b072fc8345436b7377738d53834376736a735f635a63525355535863575364636c73747375736e73757388538fd380c33a82d05260622062004200425052b8830243367359637173757382c3606342431e630e53105316531a631653165328733e834c5352535553676385c38f5383434c52f472804200422062b073024338835a6370737d837f83727368733072f472d452c442c042d052d452d052e062f8830c531a6322632e734b53737385c382c36a7343430a52e0630243434362637773844389538a53864377735e631a62c442804260624042707270728042a062c442d452f07306430e533a83687384c389d3885380c371736c73757381c3864388538743854389d388d382c37b834c52ec724041c0420042004200420042404260628852c442e8730c534853757388d38cd390d39253935393d393538fd38e538ed38a53814385c3895388d37c83747354531e62cc5220600000000000000002004200427072e4633473656384438853844387438f5392d3935393d39553965394538e5388d387438a538bd35b636c7380437e835f633272fc82c4429052707250527072b073044349537883895387437f8382438bd390d390538e538d538bd3895386c384c381c388d38e5363635d63707381c382c380436f7364635453367326633e8344434c536c7385c38cd38bd3885387c385c3824376736163515349534a534e5351535753717384436c73505340434043485359637573864387c380c37c838143824383c38b538b538ad38b5388d37b8359633e831862f882e062cc52cc52d862e8730443206343436f734c530a52b882a872d053186343435d637883844387c389d38bd38e538b538b5388d3798349530a52d052b0729862707250524042606280429862a872d0537f836873454304429052404250528852cc531c635a6376737f838143854386c38b5386435f630a52a062a062a87288524042206220622062505240426062c0437273788373735d633672f882c852905260629862f47328734c53626372737b83874386c36a733072d862a87298627072004200420042206250528852d8631e63495367637983804378835a63464332731c630442b882a8730243424365637b8386438bd38b537d8346430a52d862a0628852a062e0630243004322634d53697310534b536f738343854382437f837b83747364634b53404332733a835863788382c38543895387c37a836c7358634143434346435963697365636b737273747322634c536b7381c3874388538a5389d388d38a538d538b5382c37173687373737a837b837983767372737473717365635d63565354535653586356534e53485359636d737b8382c3874388d385c378836c7372737f8385c389d387c380c37c83788377737373636346432c731a630642ec72e062d452d052e062f472f072e8737e83824385438643874386c373734a53165300430a53206340434853434343434743535361635f6343430c52c8526062505250522062004240428042885280438bd3895386c385c3854383c36f734342f472b882a87298628852804280428852a872e46322634b53505344431a62d45288524041c041c041c04200422062206;
        // label:4
        // input_ANN = 16384'h350537a8387c388d383436563555354534f533a832063105322634643565355534343226314531c6341435c637a838c53925394d398639be39ae396d385435c6360637e8386c384436a732c730c531c6343435e635e63444332734b5360634f5328730042d452c852d4530043414373738a538f5392d39753996398638bd36a737773834383c37a8367634b53206308532c7362638243798366636b737f8370734c531252d862c042b072d453165350537b8388d38dd392d3986396d38d53747382c3854384c380437a8375735353347345436b738643895386c38743895388d37d8357531e62e462c852e0631a635153767387438e53945399e397538dd37883885389d387c381c3727360635353515360637d838b538f538e538b5389538b538dd3824351531862fc82e8730a534a5370738543905397d398e395538cd37b8387c38a5388d381436563424328733673545376738a5390538ed38ad387c38443864383436a734b53444344434743575368736f73798385c38dd38fd38b53834384438543874382c36a734853186302431c63545381438dd38fd38ad37e836b7371737e837f8375737d83834384c38343757350533a8350537c838dd3935391d364636b73767379836f735c6336730442f47320636363874388536e734b53495351535f63747387c38e53915392d38ed37f8347430643165356538543955399631a632e7341434a53565362634f5324630643165351537b8383c36a73388310530c53327366638b5392d39453955392d38ad35e631a62f4731863545382439152f47304430c5318632c73454352535053464345435e637983854380c34f530042d8631a635963844391d39863996397d394d37f834342e872f0733a8372738d5324631e6320631c6314531053327354536563697378837f83834385c373732a72dc6308534b537c838dd394d397539863986387435052f472ec73414374738d53616357534d534143287320633473586375737b837e8371736b73788381c35c6346434f536b7384438ed39353945394d393d38b536f7341431a633e836b738b53854380c37b837073626360636f73824387c383c380436463414336736063777379837473777380c388d38d538e538ed391d38fd386c3767369736d73824390538ad389d388d38853885387c38ad38e538f538bd384c3798352530c531c63606372735b633c8340435863717380c385c38b538e538cd389d3895387c38b5391d38643885389d38bd38f5391d391d38f538d538d5389d388d380c35e6336734953626354530642c442fc834853737385c38b538e538f538b537e83737381438bd388d3895389d388d386c389538c538ed38f538b538c538dd38ad383436f736973727365633072c042a8730e53555382c38f5391d38f5384435b634543575376738b5389d37f835f634a5350537073895390d38dd389d388d38853844372735d63606369735e632662c442d05341437e838e5394d3935383c34f5312531a6347438643804358631252c442ec7346437b838f53915388537f837f8380435b632063044324634e535963347312533a836b738ad394d3945385c357531252e463024388d380435052f4726062a87324636f738fd39153874377737373747356530e52b072a872fc83474368737473727376738953925393d38bd36c732e72e462dc638d5385c35b630e52a87288530a535c6388d3935392d38b537e8364634c530e52b07250529863085355537983834387438cd390d391d38ad372733672e062d0538b5387c3757353532c73085334736973895392d39653945388d36b7345431452d05270727072b0730c534a537173864389d3885389d389d37f8355531e62fc83814388d38a5384c377736e737e838bd393d3955395d393538d53834365634142fc82905260627072c0431c635c63804382c36f7369737f838ad385c36d7352534f5367637773788374737d8388d391d394d3945392d391d391538dd3814363633c82ec7270727072cc5320635753767384c372734b53454377738c5392538fd2f4730e5320631c63145330735553767388538ed38fd3905391d3905386c37f8369734442f882d05300433c835e637173844383435b632463485382c395d398628853004320630e52b8829052d45326635f6383c38ed3925393d3905385c385c385c37673525341434953646378837a8381c38243737350532663575384c390d25052d05318632e731862e462b882cc531c6360638b53975398e392d387c3854388d38953844383c384c387c38ad3895382437a83737359631a631053515377730a53105320634443575353533e830c52f07330737a8394539ce39c6397538f5389d389538cd390d3915390538f538e5384c378836b7351530c52e463246356535d6366636b73707377737883727363634e534543626387c3955395d391538ad380c372737473804389d38ed38ed38d5387c37a83717366633072e0630853444367637073747376737c83804380c37e837573676365637e838c538b5376735b6344432a7332735053767387438a5389d3895381437b837d8368731e62e0630c5359635f63646369736e737573777376736c7354533e834c536e73824375734142f072c442e8732e73636384438c538c538b5385c381c3854389535e63165300435963596352534b53495355536763717366634342f472c85300433c835c634442fc82a062c853226364638a53955393d392d38cd386c386c38cd3844361634f534b53495330730a530043165347435f63636351532872f072a872a062f8831e631452ec72e0633073777392539863955394538ed38ad389d388d3874381c380c;
        // label:0
        // input_ANN = 16384'h38a5396539a6386c36d739f6389536c7383439b63915385437b837f838ad390538443854399639a6382c360636e7387435b6354536b7384c390538fd38ed38fd3777397d399636e73424394d3a46398e38dd391d399e385436f737d8389d380c35b6367638b5382c38c5382c36873727386c37d835b63586380438ad38ed390530a536c7386c36b735153854392d3717356538b5395d38c5382437983727385c388d37c8354532a7376736c73226310535a638243834366634c5365637c8387c2d453646397539ce388d353537c838343687365637373707376737a8364635f63707382437f83606380c387c37d83656350533c834f536973626368735353586351538b53aa73b1f39fe36f73864395d386435753676387c391d38bd3814381c387438f538a53535351535e636e7385c38dd34f531a63485360637b835e6342439d6393d393d3a263a7e385437f83844384437a83717388d38fd390d39ee395536b735a637c836f735f631862f47360638c53895381c368732c73464359634c53a7e374735e638b539a636f736a7364635253515360635a6340433a83666362633e8352538743804382c3727355534a534d5375737c8364635f63606343431453a5e36a73545383c397d38ed37f836263616382438ad372734a53367340436a7385438543636316536a7399638ed347433a8330730a532063757384c363634043a56390d3844381c380c387c38cd38fd39963a873a2639a6395d392538ed395d39fe391535b63414386c3a0e39753844388d355533e836d738b536a734b53555389d38a538cd37e834a535a6389d39a6396d389d383c392d39c6397538f537e8380c38b5391538fd39c6388d366638243a06398e38743844382432c72c4430c536563707382c380435f6361635f63656362634b53474352535c63596345430a5308535f638e5373737a8346431253717398e39ce3905387c3844348532873266368737d8379837f838743525312531a63555380437e835b635353606357534c53535380c38d535553737358634c538cd39b639e6398e394d3975389d37c836c73824389d38ed399639be3656355535f638343a463a0e395d38fd39153965399e399e3986393d38e5397d397d39453915376738c53814361638a5372734a535a638bd38853915397d390d3895394d39d639c638fd3656370736e7366638d5398e388535a63515391d3a0e3a8f39b63646324634f533673246382434f533883606386c364637573767359638dd39ae38ad36f735c630c5338834343226347435d6358633a8336737673788392d39863656351535e634d535a63986380435c63565380c356537d8385c3535364638b536d733c8360635c637d83864374735c635f637f8388d37c834b531e637a839fe3945396d39c639a639c63a2e36d73505355538ed37a836f7381c37c8324636d738a538ad39553975398639ae39be39863965397539c6392d353534953707380c376739be3acf3a6e39ae391d36a7382c396538f53727353537d839a636c73747392539de394d38fd3757372738ed39f639b6386c371737c83915390d36973307354539ae397d3854388d39f639d63a2e39e6382437e8372738743a5e3a1e3834364635a634f5352531253388382438853505359637d8389d3a0e3a1637b834e53798391d34e5343438ed3a66380c38643925380c399e39ce393d39a63aaf387c348531e63307352533a835e638c536e72f4735253945397d3874390d390d3905399e38d534a5364639ae38cd3307368739de381c39ae39fe382c35e6399e39ae386c374737f838d53874386c38ed386c3515382c393d3626318636d73915396d397d399e3915397d39d6386c36a739053a76365637f8394d37d832c7387439a6399e3935390d398e38ad35f635f6398638dd38ed38a535b631c6380c38cd36e73646395d39fe39b639b63a2e39ce38f538d53404354538e539053636381c3616362636f735e638c538b536e737883a1e383435c637e83975387c39c63824332734f538fd37b8368738ed3a5638643545369735d63737394d3a4e39b6388d336731e63388320638953a0e39c63945393537d8371738d53a6e39d63935386c382c38a5384432e73434389d38e536e737e838f538bd37d8379838e539de396d3757359635153474368738cd38bd3646347438a5397d386c36b736f73616389d3a3639ae38cd3814386c383c3575388d38b538543945354530e533a837673a0e39fe390d3874377732263535360632263105390d38c533882ec73656383c37f837d838cd3a0639f6390d383c381c385c35f63606391535f633a8344435b6389d393d38f538ed38dd34343616380436c736c739de384c3287338838e5389d342432a7384c387c35753606394d3a87390d389d389d390538dd38ed38cd36d733473697389d392d399638e5395d3a1e39ce388d389d390538dd38c539be386c35e63737392535053145350538ad3a063abf3a26383c397d39c63a5639e636d730243626388d38dd39be39be397538e5380c364635e63925399e37d838dd39de39ae393538fd380c363634e53646397d3a8f3a4e399639ae39b63a4e3a16385c3656375735b634d5376735c6360635b6361638d5392d38dd35e63226386c391d388d37073646392d386c370736f7374739153a2639b63636388d3a2e3abf3a763a26384433a8314534a530a535f638d538fd38d5396538d5375736873747343435b63844382c397539ee388d35d63687392537d834443004368739b639ee391d3a1639253687359637d836a7391d39c637673246363638bd3996393d361634f536f7375735b639153a8f39b638d539f63a0e38243727;

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv1_hex.txt", "r");
        for (i = 0; i < 6; i = i + 1) begin
            code = $fscanf(fd, "%h", memory1[i]);
        end
        for (i = 0; i < 6; i = i + 1) begin
            Conv1F[i*5*5*16+:5*5*16] = memory1[i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv2_hex.txt", "r");
        for (i = 0; i < 16; i = i + 1) begin
            code = $fscanf(fd, "%h", memory2[i]);
        end
        for (i = 0; i < 16; i = i + 1) begin
            Conv2F[i*5*5*6*16+:5*5*6*16] = memory2[i];
        end

        fd = $fopen("D:/Material/CSDP/Data/Weight/distilled/conv3_hex.txt", "r");
        for (i = 0; i < 32; i = i + 1) begin
            code = $fscanf(fd, "%h", memory3[i]);
        end
        for (i = 0; i < 32; i = i + 1) begin
            Conv3F[i*3*3*16*16+:3*3*16*16] = memory3[i];
        end



        fd = $fopen("D:/Material/CSDP/Data/small_test_image.txt", "r");
        for (i = 0; i < 10000; i = i + 1) begin
            #(PERIOD / 2) reset = 1'b0;
            #(PERIOD / 2);
            status = $fscanf(fd, "%h", input_ANN);
            #((75050 + 20 + 550) * PERIOD)
            #(PERIOD * 100)
            #(PERIOD / 2)
            reset = 1'b1;
            #(PERIOD / 2);
        end
        $stop;

    end

    Lenet UUT (
        .clk        (clk),
        .reset      (reset),
        .CNNinput   (input_ANN),
        .Conv1F     (Conv1F),
        .Conv2F     (Conv2F),
        .Conv3F     (Conv3F),
        .LeNetoutput(output_ANN)
    );

endmodule
