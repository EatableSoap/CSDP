// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\IEEE162IEEE32.v
// `timescale 100 ns / 10 ps

module IEEE162IEEE32_TB ();
endmodule