// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\layer.v
// `timescale 100 ns / 10 ps

module layer_TB();

parameter DATA_WIDTH = 32;
parameter INPUT_NODES = 100;
parameter OUTPUT_NODES = 32;

reg clk, reset;
reg [DATA_WIDTH*INPUT_NODES-1:0] input_fc;
wire [DATA_WIDTH*OUTPUT_NODES-1:0] weights;
wire [DATA_WIDTH*OUTPUT_NODES-1:0] output_fc;

reg [7:0] address;

localparam PERIOD = 100;

always
	#(PERIOD/2) clk = ~clk;

layer #(
    .DATA_WIDTH(DATA_WIDTH),
    .INPUT_NODES(INPUT_NODES),
    .OUTPUT_NODES(OUTPUT_NODES)
)
UUT
(
	.clk(clk),
	.reset(reset),
	.input_fc(input_fc),
	.weights(weights),
	.output_fc(output_fc)
);

always @ (posedge clk or posedge reset) begin
	if (reset == 1'b1) begin
		address = 0;
	end else begin
		address = address + 1;
	end
end

weightMemory WM 
(
	.clk(clk),
	.address(address),
	.weights(weights)
);

initial begin
	#0
	clk = 1'b0;
	reset = 1'b1;
    // input_fc = 32*100 = 3200 bits
	input_fc = 3200'b00111110110101101010010110110100001111110011010001110101011100000011111100101101101110010110001000111110101011101000010101010100001111110110000001111111101110100011111011000011010010010111101000111111011111001000101111111100001111110111001000101111111000000011111101011010001000111010111000111111011101000000011111101110001111100010111111011001011101100011111100000010101100110000001000111110101010010111100101011010001111101100110010000101101000000011111101111011101001111111110000111110011010111101000111101110001111110110011010000011110100100011111101101111110100011101110000111110101011011010100101100100001111100001000110100001000100100011111100010001101100110010100000111111001011100010000101100100001111110111100011001101111010100011111010100100100001010011110000111111010011010100111110011100001111110010101001000011010101100011111101111100000000000000000000111110101010001011100101010110001111110100110001101111100111000011111000001100010010010011010000111111000110110111111100111000001111011001010011100001001010100011111100001100000001110001010000111111000000111101100100000010001111110110111100001011111000000011111100111000110101110110101000111111001011110010100101011110001111110110111101110111111000100011111101101001101000011100101000111111010110110100010110111110001111110011000111010101010111100011111101001000000100011001000000111110110001001110100110000000001111101111011010111101111101000011111011110100011110011111011000111101110110011001000110111100001111101110000100001101101111100011110110101010011000010101101000111111010100001000110110100000001111101011010011101101011100000011111101100000101000011011111000111110101110111001010110000000001111110100010100110011100011100011111010010001011000010001110000111101010111101000000110110000001111110101100010001101101100000011111100001101101010010010001000111111000000111001100100001010001111110110010011011011110011100011111101101111001100111101101000111111010111111011100110111110001111110001000111101011001000000011111010110001110010010111000000111111001100001010001101100010001111101010011010010001010000100011111101011110000100111100001000111101101000101100000101000110001111110110000011111011110010100011111101010010101000111010110000111111000001010101101100000010001111110010101100000101010100100011111100000001111101010000011000111111001000010011100101000010001111101100011100001101100001000011110110111001100100010111100000111110111101111001110111110100001110110111000000000001110110100011111010000110000011010000001000111111010010010011011110001110001111110000111010110101000111000011111101111101111010111111101000111111000110011001101100101100001111011000101110000001000101000011111001010010100010011001100000111110110100011001010110101010001111110011100101111011011101000011111000110011010110010111100000111111000110111101100100110100001111110000011101111011000001100011111101011111000000111100000000111111001110111111111101111010001111101100001101100101100010000011111100000100011111010000101000111100001100111000000100110110001111110110110010100011110101100011111001011000011110011100010000111110000100101010000100110000001111110101100001110101101101000011110111101101011100011111001000111101011101111110000111101110;

	#PERIOD
	reset = 1'b0;
	

	#(102*PERIOD)
	$stop;
end

endmodule