// CNN_FGPA\CNN_FPGA.sim\sources_1\new\convLayerMulti.v
`timescale 1 ns / 1 ps

module convLayerMulti_TB();

parameter DATA_WIDTH = 16;
parameter D = 1;  //Depth of image and filter
parameter H = 32;  //Height of image
parameter W = 32;  //Width of image
parameter F = 5;  //Size of filter
parameter K = 6;  //Number of filters applied
parameter P = 2;  //Number of padding pixels

reg clk, reset;
reg [0:D*H*W*DATA_WIDTH-1] image;
reg [0:K*D*F*F*DATA_WIDTH-1] filters;
wire [0:K*(H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH-1] outputConv;

localparam PERIOD = 4;

integer i,j,k;

always
	#(PERIOD/2) clk = ~clk;

convLayerMulti #(
    .DATA_WIDTH(DATA_WIDTH),
    .D(D),
    .H(H),
    .W(W),
    .F(F),
    .K(K),
    .P(P)
)
UUT 
(
	.clk(clk),
	.reset(reset),
	.image(image),
	.filters(filters),
	.outputConv(outputConv)
);
	
initial begin 
	#0
	clk = 1'b0;
	reset = 1'b1;
	#1
	reset = 1'b0;
	// input image = 1*32*32*16 = 16384 bit
	// expected output = 6*32*32*16 = 98304 bit
	 image = 16384'h33883525368736f735e633272f472c04298628042a872c852d862e87300431a633a834e53586358634d534743404324630642ec72ec730e534143606377737673676370737a837d83727351531652c4425052004200424042505260629052c442f47314533273454341434443505359634e5332730e52f472f88310532a73414377737983777379837e83788359631862a87240422062606270724042004240428852c442fc8326634443575367636c7368736c736d7362634c531a62f072e4636d73656366636f737c8385c3854369733882ec72a062707240420041c041c04200427072cc530c5342435e6363634e53307342435653666371736b735d634f536c736763717381c386c387438b5388d3788355532e72fc82b88288525052206240428852d053186350536b73697347430642e062f073165348536c7380c380437c8385c387c38b538fd38d538a538ad38b53864379835a633e831e630c52fc83004302430e533e8365637a837a836a73505338831e6318632c73535372737f8388d390538d53874383c37c83798384438d538fd38dd3854379836d7363635b635e63616363636d737f8384c383437c837073505324630a531e634a536873767390d391d388536d73485324632e735653788386438d538bd388d3874386c3834385c388d388d388538a538a5386c380c371734442f472a062c043044347435f6395d3925383c354530442b882c042f8832e735a6381438b538cd38c538d538ad389538ad38dd38c538dd387c381c37e8371734c531c62f472c042986306434443975396538c5363630852a0629052b072dc631e63616384c38c538cd38ed38d53895389538a5383437983656353534d5354535453555351533e8310531e63474399e39ce392d37c834c530042c442cc52e873125352537c8389538dd392d391538d538dd387435d6334731252fc82e873044320634743616371736c7369736b7399e39ae3965390d38543565338833a8347434d53626380c38b538ed38ed38ed38f538cd37a833a82ec72c042986280429862cc5304433883646381c3854380c397d394d394d3986396538a53824380c3814380c3834387438ad388d3814382438a53874363631a62cc5290526062206240428042a062dc6328735c6377737b8392d38c538d5390538ed38a5384c3834382c382c38743885386c380c37073737385c388536c732462c442707240420042004240427072b072fc8345436b7377738d53834376736a735f635a63525355535863575364636c73747375736e73757388538fd380c33a82d05260622062004200425052b8830243367359637173757382c3606342431e630e53105316531a631653165328733e834c5352535553676385c38f5383434c52f472804200422062b073024338835a6370737d837f83727368733072f472d452c442c042d052d452d052e062f8830c531a6322632e734b53737385c382c36a7343430a52e0630243434362637773844389538a53864377735e631a62c442804260624042707270728042a062c442d452f07306430e533a83687384c389d3885380c371736c73757381c3864388538743854389d388d382c37b834c52ec724041c0420042004200420042404260628852c442e8730c534853757388d38cd390d39253935393d393538fd38e538ed38a53814385c3895388d37c83747354531e62cc5220600000000000000002004200427072e4633473656384438853844387438f5392d3935393d39553965394538e5388d387438a538bd35b636c7380437e835f633272fc82c4429052707250527072b073044349537883895387437f8382438bd390d390538e538d538bd3895386c384c381c388d38e5363635d63707381c382c380436f7364635453367326633e8344434c536c7385c38cd38bd3885387c385c3824376736163515349534a534e5351535753717384436c73505340434043485359637573864387c380c37c838143824383c38b538b538ad38b5388d37b8359633e831862f882e062cc52cc52d862e8730443206343436f734c530a52b882a872d053186343435d637883844387c389d38bd38e538b538b5388d3798349530a52d052b0729862707250524042606280429862a872d0537f836873454304429052404250528852cc531c635a6376737f838143854386c38b5386435f630a52a062a062a87288524042206220622062505240426062c0437273788373735d633672f882c852905260629862f47328734c53626372737b83874386c36a733072d862a87298627072004200420042206250528852d8631e63495367637983804378835a63464332731c630442b882a8730243424365637b8386438bd38b537d8346430a52d862a0628852a062e0630243004322634d53697310534b536f738343854382437f837b83747364634b53404332733a835863788382c38543895387c37a836c7358634143434346435963697365636b737273747322634c536b7381c3874388538a5389d388d38a538d538b5382c37173687373737a837b837983767372737473717365635d63565354535653586356534e53485359636d737b8382c3874388d385c378836c7372737f8385c389d387c380c37c83788377737373636346432c731a630642ec72e062d452d052e062f472f072e8737e83824385438643874386c373734a53165300430a53206340434853434343434743535361635f6343430c52c8526062505250522062004240428042885280438bd3895386c385c3854383c36f734342f472b882a87298628852804280428852a872e46322634b53505344431a62d45288524041c041c041c04200422062206;
     // filters = 6*1*5*5*16 = 2400 bit
	 filters[0*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h9820b02b2c172bddae3120351d7e2a55b4f1313c2dbd2b5f33c631b1248d28162fb2a9c4a6c932d3175bb01fb374a549b125;
  	 filters[1*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'hae582e0dabad2c8a28e42af1a0662ea42fe0a6629a3faef3b912b05b2321339a3067b83ba2f12cd12fd335a0279630cea62e;
	 filters[2*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'hb680ae8c2a85a7322b32b66833c8350732102d2ab15a35742ae5b4f9afa0307e29359e1eaccb2ecc2f24b051a0072ce6ab5a;
	 filters[3*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h29e5220c33e6b287aac2286f356e3198b210afc32b4930db2fc8b5a0b29026c0274427e5ac67ae352ea1ac83b00e2a622498;
	 filters[4*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h2bc0af8f31742da42f32b0d631e131aa347631442dc7ad87a44cb231ac5e2d2f247bb4b5b7eda68e2b7aa8d99fd5ac7fad33;
	 filters[5*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 400'h31e1b46a2dce34d4acb8ad1eb6ff30be374e2aa931e0b6a1a538aca02cd9b0942f6eb12da9b628b71e8a9c7ba5d02e70a93b;
	#(PERIOD)

	// reset = 0;
	
	#(3*1793*PERIOD)
	// Display output
    for (k = 0; k < 6; k = k + 1) begin
        $display("Kernel %d result is %h ", k+1, outputConv[k*(H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH +: (H-F+1+2*P)*(W-F+1+2*P)*DATA_WIDTH]);
        $display("\n");
    end
	$stop;
end

endmodule
