// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\UsingTheRelu.v
`timescale 1 ns / 10 ps

module UsingTheRelu_TB ();
endmodule
