// CNN_FGPA\CNN_FPGA.sim\sources_1\imports\Integration first part\convLayerSingle.v
`timescale 1 ns / 1 ps

module convLayerSingle_TB ();

parameter DATA_WIDTH = 16;
parameter D = 1;  //Depth of the filter
parameter H = 32;  //Height of the image
parameter W = 32;  //Width of the image
parameter F = 5;  //Size of the filter

// tag: convLayerSingle.v is [0:n-1]
reg clk, reset;
reg [D*H*W*DATA_WIDTH-1:0] image;
reg [D*F*F*DATA_WIDTH-1:0] filter;
wire [(H-F+1)*(W-F+1)*DATA_WIDTH-1:0] outputConv;

localparam PERIOD = 2;

integer i, clkCounter;

always
	#(PERIOD/2) clk = ~clk;

always @ (posedge clk) begin
	clkCounter = clkCounter + 1;
end

convLayerSingle #(
    .DATA_WIDTH(DATA_WIDTH),
    .D(D),
    .H(H),
    .W(W),
    .F(F)
)
UUT
(
	.clk(clk),
	.reset(reset),
	.image(image),
	.filter(filter),
	.outputConv(outputConv)
);

initial begin
	#0
	clkCounter = 0;
	clk = 1'b0;
	reset = 1;
	// LeNet first layer = 1*32*32*16 = 16384 bit
	image = 16384'h3971328133ed36953a0a250f3594380933e5357239b827103009375e36fc375638932d04323635e9388b394a35af3b87378e359d31fe376f387035db35f6332a3a64384036bc3458387539db351b366838a83808302b3742395e3764382c38a73ac934333a823a0438c83b6e3a6639893ba83b9837bb393433a127ab270335ac3a933985369839023aaa32fc3650319d3a3636c2345932a530da31e91f9034d7383d30fc387c36893a963480395d3a33362c30eb35e73707332b33af372d25633bf0377d26b0367b39a1341939db3b8a3250212f3b4c352038e4349832a733ee34283a352cdc379b3af4353538b93a6138da34c13b8f38093bd636de38a33a68349a24a73bb43ba03489398e2626388438f838142b5f222138693ad03b3c38253a12383e271836502ec638b234593b9039ce368a336738a6389d35ab38503a9b382d2eed317b348e3af232202c553a5c3b1236ed3beb38a031dd388a3ac53b5b36dd382d2ff239b936763a3434e833d536fd37f13ba136e139a63abb383c253b38483b2430503b1d38da32bf34b5340834a2396539661d303afb3aab39753b6138a035ac3bf2380322ad3a61393f345f389e2c9132353a9b38ca3a47339338dc382335b134ab3851365339f2385039c43b6537b0390238023ab829d3399a36f9389f39b13be136933b58391639e73b383762399739a2308938f537dd3a52344f30b03a432fc339203b2c2f303aa636832a5838cb38493bf8392135b6343e3b0b37933833334239dd3b0c3bdf395133ab3ab738d732b0302d3941380236403bba3680393d3b4221d4316a3aa13bfe23f81bcf31ce38d73777275b31d72a112c22399d398737242fdb37d4381d369f39aa2613394438d93abd380e36a534843b07387f38b4382032823b123189356232c630393aca3377385d343a32272ede34023433383e381639ff39e13883349b34bd2eb438c637a53415363a36742a48393e37a23bc43ac832ef33f737aa2d3633e6380338b032b93324359c31513014394430753b9237a73a1538022e2a31253a1d393e3b1c358538373030396924861ecb22373a0d3bda3aa72eea3bff37903b88362734bd395736af39e539d82022393539f13b963ad739293a4b331b3a1139793b283239391a3bf82b39361c3ab73b2838f23abf322a395135593bc9358d36d03b9128fa388d39ba3b8b39f239643574395d3afc374438e73bac1fbc36cd379f36113838359c30812db13595364039c73b6a319338fb35ac301d2d133a8d2000307d39b939242d7138ba3b2d3992377339ef3a84341f39cc39bc35d53a72340632753a5131ec34b4381b36e93a862eee32703be138af35fa360335b43a5f35ee34ba3088300c3715380638323a45354f3ad737c2391f3b131cb33278323635563a633ab834063489362232aa3414397f3549349739c62dc72ea437e53b5b35603b9d387938b42af035ab36f73a2535ce3341388b2763388736c934663b40302d3b4d33563a5d390d336b3bf6366a39be37da24f93599254937142ff63814341836af2ee2394826c73b0b301b365a35302a91395e32753b5e32ec3ba938e53a2d3b2c3b8c39ea35263b753b3c3b5a2f29333c38e43a172e9234f33b21394930e438ab380033db35183ae73a6d39e02f2e3bfb2d6b38fc374e377e38be35673a7c3008265b35cd344c1990355137ee383b36af26293b9c385f36c731bf386b3950375d30e63bbc3a63379c38be34f3350a35a63a0c39733aca3965397d3a813bfd3b9232eb3a143aee388d39e238d52bda3bea383038c939722b2034e22c2a39f536213854395a394e37943b6d3afa378a30ea3986398339643749399938b03b213b2e33013b9536c934e7320334b93639382c3bfe354833ff300c3a48373f3bb931d026f53b2f2a4431b73a3b31fe335738cb37f230df393e39e83abf3bc23ac239db230f3906309c3bfc33b33a35382b36c9319738163ab833c9296435b839a334e338ae37aa289f185438b537d33ba33b1e3a94340b3b8638733ad63287356d3b8e2123375b36753539372d36ca37843604397c2646336335593bde3a1e32f935d434de3bd4394339bf379330c73b372a483b3e363f3a6b3b48392336573b8a3a6436183b5b3a043af139ab3a753244302335a6385a370231683a11382c27a93ac4388d3083393d35cc2dc43a792f5835763b28376738ff3aaa393638993b0d3a2b39ca399034ea353d3bfd24653ad136f23b843117366e2e953bd238e234043aa13aeb38bd3b3638943b28395939b129c124f638f3374234bd389834643b7c32833b3d3beb3aa035722a3a32d735da373630f5310038832e5738df32703a263b2e3a1f372438af361038fc3b432fce33d839ca357b31983bf836c02fbe2f1a3add3a4338b73b203ad13a7b37cc381f381137ad3ac0331839cb37d73ad628d539393964385c35643a0239f03bff38f1379430143854356b3a5b2d3c39b83a8637e73baf36bc329c38fd388338b43a3737a030e3360f328b3ad33a0237d73585398e3a9238923919304e35933a5838023ac73b853abe34b03b34386a39b03a9633673a0a3781379138c338d5355439793af4388f39e13a0e34a53b613bed3bec39273a3d31472e61395737f9374239462a823a4b38cc3ae63b1937ac39e43880341d3bd433bd36312deb366f390032803776333b3a103bcc394a26212ca93a6d38f6301c2e5635cc33f32fbf39f7396a3663310a2c03386d31ba3b9534f33b1a3515396b35792f003a833b37369f369b3bf0317b2fe73bab38023816380b31ab39e834de38652f3731493a9a30c932b038dd32c738c335bc3aca30fa39f83b2e339a3254334b38c539fa386e3bcf39b8;

    // filter = 1*5*5*16 = 400 bit
	filter = 400'h32fd248a377eb43cb630b3d6b31335de35702dadab7c37fcb6b3b6c7b707b336ad61b411b7e1b71b33473523b65d35fc379c;

	#PERIOD
	reset = 0;

	#((56*28+1)*PERIOD)
	// for (i = 28*28-1; i >=0; i = i - 1) begin
        // $display("Result (hex): %h", outputConv[i*16+:16]);
	// end
	$display("Result (hex):%h",outputConv);
    if(outputConv == 12544'h55585d7e5b9759f25d375582548f5f865e3c584255485da95586574655ab5d6a5c8258c25b5c55635c0c5a74cfbe5f8d593e5e1957d455ff57ee5ea053725bf35a7c56175a965c5a5de0592a5ada561b5cad58765bf056005ab25c7157d0592b5966c75e59b25f135ba95e115c2c5a375be55c1b564e57225d8f5a805d8258775d5e59055a535698d3065e695c165dd95875591c59f65d0854f95b0559d25c7b4c745d915ba85abf5b37524a59c15c5b5828591d54905bf45ce65d7858755ba15a315d54d1bc596054675e05559957005b745bda5b0e57865b315ea558215c6558ec5ab657a9567355f35d79522359db5d1a54175e485a5451225ae95c0c5ac55c3750795c30591952785a3959d75ce651315c925bd459b8d0ea541251d15c905a19cc8a5c9d5c845dee5b04595059b45c3f51d35a0b5fbb54915bcd5b4f5a6f44d65d9159175b9e553459935b765c80583254385f03558f5cf45bcf59e45be05d16570e5963602d5bfd5c3a4cb05d8dd0365d295c2c58d258755c80566e5a085b845b35557e5b2658d15d90596c58465d195a4753695b45525a58ae5bd55cfd5a4959ec59a85e225a3b5e18580155e45ba2d77a534c5aef5d365e565c095e3f5c41595d55205da95b1f5ab3d24659de59e3597559555af35aae5ca55a46587553785d085d3d5a025b724eb959f054d058c65a2e5b3b5a6d586558e15cba59095aa35a3658405b9654975a12571a5d485a625e965ce15d6e51f15b474e54590355b35c045d1d4e785abd55eb5b8a5b935f1752cc5c17593b5cba5c0b5cbf58ba5b3b54555b325b835a745dc85b725a09d42b59dc5a205c2a58f053425dc04c875b3e54385c895e085a08582d5d2c5c885b33583d59255c9159065add5c5b59a8551459325ccd5ea7d40150f0551559935ce55cc359a057c55ae253c550895b2d58c1580758e75946587e5c3d5a255cf858025c3154975b2fce93575259ff5d424fda5dd0560a512f5a2257db59975d255b074a8b5abc5abc5f2658b65b38cea559aa5b245c425a905d3d5a5a540a575455525c395e64581fd6975ffc51ab50c45c6351a45a005a775de558a95c0858245d1257ea5e115d465b494a405ce4cf1a5bcc53615d135c605ba95ae45b81c4635abb5d4bd17359ae5e9356185f444a365b915be35a9f56175ccd55605a18558d4a7359785b86cd5f5d2556105d07597654f054f35be75bf850ef6012d01059c458794c875d665d785ca55c8358de5045588d5da85c905c8c5c3d5928595a596d585959ce58ee570254305cb54dd25a8cd4b45bb057235e425aad54f75cd0ce655bec55895be05a8e4d24405b599a5df05c115ae05c0f599d59e858115af258fb5c86beda5cc05a345bcc5c1856045aa358a754fc5b88595e58dd586858ad58bb5a8458175cf95c895dbc5aac5c7158805d0155d3d0115b7a5c17592556775ccb583b5ef456ca5ac6592e597b5b5e534e5e265561588d5b10583b58df5d0e5c7b5d63590b574c5a155cb15a4dd3695c015c055d7f5acb583959245cca5b815a345ef356be556650bb584546c05f8958bf5b8b5b8358c55abf5acd5c2644985ba556875a315c355e5f5b9359015d7d550a587b5857562654385e985b0559705c4d5675589b55f8591558ad5e2258d34c1259205a60538a5f875ba05c525a47cf7757995b835dee59635b1f5c5655cb5cc15938474956085b574daf5bac59df5b38592f5a5c5a46557f5ad95b8b5b5b5c5e581a5b075c2e58cd58645cd35990591b592f5bd1cde45c2d58de5b515d955811571fd2305cd74bc055fd5ee0594158ba5e115a5a5bcf5c35579b5c31585f5a395ca753cd59c25d085dc556a5d424590e5c0ed2485bef571c5ea9589959a54e2f598b5ef35cb65c825cb9d4b352875b3e56175d205cba57085f4d3fd359b558f65ac2570158525e1a57615c385c1bcc4359b858be56285ddc59f55cac4a465d1e5a53580459145d1bcc4058d75ab9587c5dd756505d46550f572e5b025d7c59e357fb5ab65aed5c135bee5c40584f570b591156f0599458ae5ba75b415d2f54ed529b5cff5a9a5b215b485bdb5d4855ad5ca159b758f559ff54355e82571851945cbd5bb959f85c78588255314d285f105a055aa85c4859afcc85559f4ffc5c9e5e4a5b645e13cabd5a73553e5903593e5a0354425d3a5c645a5fcaf25c605dfa)
        $display("TEST PASSED!");
    else
        $display("TEST FAILED!");
	$stop;
end

endmodule